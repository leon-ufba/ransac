// RANSAC_NIOS.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module RANSAC_NIOS (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] processador_data_master_readdata;                            // mm_interconnect_0:Processador_data_master_readdata -> Processador:d_readdata
	wire         processador_data_master_waitrequest;                         // mm_interconnect_0:Processador_data_master_waitrequest -> Processador:d_waitrequest
	wire         processador_data_master_debugaccess;                         // Processador:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:Processador_data_master_debugaccess
	wire  [18:0] processador_data_master_address;                             // Processador:d_address -> mm_interconnect_0:Processador_data_master_address
	wire   [3:0] processador_data_master_byteenable;                          // Processador:d_byteenable -> mm_interconnect_0:Processador_data_master_byteenable
	wire         processador_data_master_read;                                // Processador:d_read -> mm_interconnect_0:Processador_data_master_read
	wire         processador_data_master_write;                               // Processador:d_write -> mm_interconnect_0:Processador_data_master_write
	wire  [31:0] processador_data_master_writedata;                           // Processador:d_writedata -> mm_interconnect_0:Processador_data_master_writedata
	wire  [31:0] processador_instruction_master_readdata;                     // mm_interconnect_0:Processador_instruction_master_readdata -> Processador:i_readdata
	wire         processador_instruction_master_waitrequest;                  // mm_interconnect_0:Processador_instruction_master_waitrequest -> Processador:i_waitrequest
	wire  [18:0] processador_instruction_master_address;                      // Processador:i_address -> mm_interconnect_0:Processador_instruction_master_address
	wire         processador_instruction_master_read;                         // Processador:i_read -> mm_interconnect_0:Processador_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;         // mm_interconnect_0:jtag_avalon_jtag_slave_chipselect -> jtag:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;           // jtag:av_readdata -> mm_interconnect_0:jtag_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;        // jtag:av_waitrequest -> mm_interconnect_0:jtag_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;            // mm_interconnect_0:jtag_avalon_jtag_slave_address -> jtag:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;               // mm_interconnect_0:jtag_avalon_jtag_slave_read -> jtag:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;              // mm_interconnect_0:jtag_avalon_jtag_slave_write -> jtag:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;          // mm_interconnect_0:jtag_avalon_jtag_slave_writedata -> jtag:av_writedata
	wire  [31:0] mm_interconnect_0_processador_jtag_debug_module_readdata;    // Processador:jtag_debug_module_readdata -> mm_interconnect_0:Processador_jtag_debug_module_readdata
	wire         mm_interconnect_0_processador_jtag_debug_module_waitrequest; // Processador:jtag_debug_module_waitrequest -> mm_interconnect_0:Processador_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_processador_jtag_debug_module_debugaccess; // mm_interconnect_0:Processador_jtag_debug_module_debugaccess -> Processador:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_processador_jtag_debug_module_address;     // mm_interconnect_0:Processador_jtag_debug_module_address -> Processador:jtag_debug_module_address
	wire         mm_interconnect_0_processador_jtag_debug_module_read;        // mm_interconnect_0:Processador_jtag_debug_module_read -> Processador:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_processador_jtag_debug_module_byteenable;  // mm_interconnect_0:Processador_jtag_debug_module_byteenable -> Processador:jtag_debug_module_byteenable
	wire         mm_interconnect_0_processador_jtag_debug_module_write;       // mm_interconnect_0:Processador_jtag_debug_module_write -> Processador:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_processador_jtag_debug_module_writedata;   // mm_interconnect_0:Processador_jtag_debug_module_writedata -> Processador:jtag_debug_module_writedata
	wire         mm_interconnect_0_memoria_s1_chipselect;                     // mm_interconnect_0:memoria_s1_chipselect -> memoria:chipselect
	wire  [31:0] mm_interconnect_0_memoria_s1_readdata;                       // memoria:readdata -> mm_interconnect_0:memoria_s1_readdata
	wire  [15:0] mm_interconnect_0_memoria_s1_address;                        // mm_interconnect_0:memoria_s1_address -> memoria:address
	wire   [3:0] mm_interconnect_0_memoria_s1_byteenable;                     // mm_interconnect_0:memoria_s1_byteenable -> memoria:byteenable
	wire         mm_interconnect_0_memoria_s1_write;                          // mm_interconnect_0:memoria_s1_write -> memoria:write
	wire  [31:0] mm_interconnect_0_memoria_s1_writedata;                      // mm_interconnect_0:memoria_s1_writedata -> memoria:writedata
	wire         mm_interconnect_0_memoria_s1_clken;                          // mm_interconnect_0:memoria_s1_clken -> memoria:clken
	wire         mm_interconnect_0_memoria_dados_s1_chipselect;               // mm_interconnect_0:memoria_dados_s1_chipselect -> memoria_dados:chipselect
	wire  [31:0] mm_interconnect_0_memoria_dados_s1_readdata;                 // memoria_dados:readdata -> mm_interconnect_0:memoria_dados_s1_readdata
	wire         mm_interconnect_0_memoria_dados_s1_debugaccess;              // mm_interconnect_0:memoria_dados_s1_debugaccess -> memoria_dados:debugaccess
	wire  [13:0] mm_interconnect_0_memoria_dados_s1_address;                  // mm_interconnect_0:memoria_dados_s1_address -> memoria_dados:address
	wire   [3:0] mm_interconnect_0_memoria_dados_s1_byteenable;               // mm_interconnect_0:memoria_dados_s1_byteenable -> memoria_dados:byteenable
	wire         mm_interconnect_0_memoria_dados_s1_write;                    // mm_interconnect_0:memoria_dados_s1_write -> memoria_dados:write
	wire  [31:0] mm_interconnect_0_memoria_dados_s1_writedata;                // mm_interconnect_0:memoria_dados_s1_writedata -> memoria_dados:writedata
	wire         mm_interconnect_0_memoria_dados_s1_clken;                    // mm_interconnect_0:memoria_dados_s1_clken -> memoria_dados:clken
	wire         irq_mapper_receiver0_irq;                                    // jtag:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] processador_d_irq_irq;                                       // irq_mapper:sender_irq -> Processador:d_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Processador:reset_n, irq_mapper:reset, jtag:rst_n, mm_interconnect_0:Processador_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [Processador:reset_req, rst_translator:reset_req_in]
	wire         processador_jtag_debug_module_reset_reset;                   // Processador:jtag_debug_module_resetrequest -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [memoria:reset, memoria_dados:reset, mm_interconnect_0:memoria_reset1_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [memoria:reset_req, memoria_dados:reset_req]

	RANSAC_NIOS_Processador processador (
		.clk                                   (clk_clk),                                                     //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                             //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                          //                          .reset_req
		.d_address                             (processador_data_master_address),                             //               data_master.address
		.d_byteenable                          (processador_data_master_byteenable),                          //                          .byteenable
		.d_read                                (processador_data_master_read),                                //                          .read
		.d_readdata                            (processador_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (processador_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (processador_data_master_write),                               //                          .write
		.d_writedata                           (processador_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (processador_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (processador_instruction_master_address),                      //        instruction_master.address
		.i_read                                (processador_instruction_master_read),                         //                          .read
		.i_readdata                            (processador_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (processador_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (processador_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (processador_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_processador_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_processador_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_processador_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_processador_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_processador_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_processador_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_processador_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_processador_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                             // custom_instruction_master.readra
	);

	RANSAC_NIOS_jtag jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	RANSAC_NIOS_memoria memoria (
		.clk        (clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_memoria_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoria_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoria_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoria_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoria_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoria_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoria_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                     // (terminated)
	);

	RANSAC_NIOS_memoria_dados memoria_dados (
		.clk         (clk_clk),                                        //   clk1.clk
		.address     (mm_interconnect_0_memoria_dados_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_memoria_dados_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_memoria_dados_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_memoria_dados_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_memoria_dados_s1_write),       //       .write
		.readdata    (mm_interconnect_0_memoria_dados_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_memoria_dados_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_memoria_dados_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                            // (terminated)
	);

	RANSAC_NIOS_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                   (clk_clk),                                                     //                                 clock_clk.clk
		.memoria_reset1_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                          //      memoria_reset1_reset_bridge_in_reset.reset
		.Processador_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // Processador_reset_n_reset_bridge_in_reset.reset
		.Processador_data_master_address                 (processador_data_master_address),                             //                   Processador_data_master.address
		.Processador_data_master_waitrequest             (processador_data_master_waitrequest),                         //                                          .waitrequest
		.Processador_data_master_byteenable              (processador_data_master_byteenable),                          //                                          .byteenable
		.Processador_data_master_read                    (processador_data_master_read),                                //                                          .read
		.Processador_data_master_readdata                (processador_data_master_readdata),                            //                                          .readdata
		.Processador_data_master_write                   (processador_data_master_write),                               //                                          .write
		.Processador_data_master_writedata               (processador_data_master_writedata),                           //                                          .writedata
		.Processador_data_master_debugaccess             (processador_data_master_debugaccess),                         //                                          .debugaccess
		.Processador_instruction_master_address          (processador_instruction_master_address),                      //            Processador_instruction_master.address
		.Processador_instruction_master_waitrequest      (processador_instruction_master_waitrequest),                  //                                          .waitrequest
		.Processador_instruction_master_read             (processador_instruction_master_read),                         //                                          .read
		.Processador_instruction_master_readdata         (processador_instruction_master_readdata),                     //                                          .readdata
		.jtag_avalon_jtag_slave_address                  (mm_interconnect_0_jtag_avalon_jtag_slave_address),            //                    jtag_avalon_jtag_slave.address
		.jtag_avalon_jtag_slave_write                    (mm_interconnect_0_jtag_avalon_jtag_slave_write),              //                                          .write
		.jtag_avalon_jtag_slave_read                     (mm_interconnect_0_jtag_avalon_jtag_slave_read),               //                                          .read
		.jtag_avalon_jtag_slave_readdata                 (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),           //                                          .readdata
		.jtag_avalon_jtag_slave_writedata                (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),          //                                          .writedata
		.jtag_avalon_jtag_slave_waitrequest              (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),        //                                          .waitrequest
		.jtag_avalon_jtag_slave_chipselect               (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),         //                                          .chipselect
		.memoria_s1_address                              (mm_interconnect_0_memoria_s1_address),                        //                                memoria_s1.address
		.memoria_s1_write                                (mm_interconnect_0_memoria_s1_write),                          //                                          .write
		.memoria_s1_readdata                             (mm_interconnect_0_memoria_s1_readdata),                       //                                          .readdata
		.memoria_s1_writedata                            (mm_interconnect_0_memoria_s1_writedata),                      //                                          .writedata
		.memoria_s1_byteenable                           (mm_interconnect_0_memoria_s1_byteenable),                     //                                          .byteenable
		.memoria_s1_chipselect                           (mm_interconnect_0_memoria_s1_chipselect),                     //                                          .chipselect
		.memoria_s1_clken                                (mm_interconnect_0_memoria_s1_clken),                          //                                          .clken
		.memoria_dados_s1_address                        (mm_interconnect_0_memoria_dados_s1_address),                  //                          memoria_dados_s1.address
		.memoria_dados_s1_write                          (mm_interconnect_0_memoria_dados_s1_write),                    //                                          .write
		.memoria_dados_s1_readdata                       (mm_interconnect_0_memoria_dados_s1_readdata),                 //                                          .readdata
		.memoria_dados_s1_writedata                      (mm_interconnect_0_memoria_dados_s1_writedata),                //                                          .writedata
		.memoria_dados_s1_byteenable                     (mm_interconnect_0_memoria_dados_s1_byteenable),               //                                          .byteenable
		.memoria_dados_s1_chipselect                     (mm_interconnect_0_memoria_dados_s1_chipselect),               //                                          .chipselect
		.memoria_dados_s1_clken                          (mm_interconnect_0_memoria_dados_s1_clken),                    //                                          .clken
		.memoria_dados_s1_debugaccess                    (mm_interconnect_0_memoria_dados_s1_debugaccess),              //                                          .debugaccess
		.Processador_jtag_debug_module_address           (mm_interconnect_0_processador_jtag_debug_module_address),     //             Processador_jtag_debug_module.address
		.Processador_jtag_debug_module_write             (mm_interconnect_0_processador_jtag_debug_module_write),       //                                          .write
		.Processador_jtag_debug_module_read              (mm_interconnect_0_processador_jtag_debug_module_read),        //                                          .read
		.Processador_jtag_debug_module_readdata          (mm_interconnect_0_processador_jtag_debug_module_readdata),    //                                          .readdata
		.Processador_jtag_debug_module_writedata         (mm_interconnect_0_processador_jtag_debug_module_writedata),   //                                          .writedata
		.Processador_jtag_debug_module_byteenable        (mm_interconnect_0_processador_jtag_debug_module_byteenable),  //                                          .byteenable
		.Processador_jtag_debug_module_waitrequest       (mm_interconnect_0_processador_jtag_debug_module_waitrequest), //                                          .waitrequest
		.Processador_jtag_debug_module_debugaccess       (mm_interconnect_0_processador_jtag_debug_module_debugaccess)  //                                          .debugaccess
	);

	RANSAC_NIOS_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (processador_d_irq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                            // reset_in0.reset
		.reset_in1      (processador_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),            // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),        //          .reset_req
		.reset_req_in0  (1'b0),                                      // (terminated)
		.reset_req_in1  (1'b0),                                      // (terminated)
		.reset_in2      (1'b0),                                      // (terminated)
		.reset_req_in2  (1'b0),                                      // (terminated)
		.reset_in3      (1'b0),                                      // (terminated)
		.reset_req_in3  (1'b0),                                      // (terminated)
		.reset_in4      (1'b0),                                      // (terminated)
		.reset_req_in4  (1'b0),                                      // (terminated)
		.reset_in5      (1'b0),                                      // (terminated)
		.reset_req_in5  (1'b0),                                      // (terminated)
		.reset_in6      (1'b0),                                      // (terminated)
		.reset_req_in6  (1'b0),                                      // (terminated)
		.reset_in7      (1'b0),                                      // (terminated)
		.reset_req_in7  (1'b0),                                      // (terminated)
		.reset_in8      (1'b0),                                      // (terminated)
		.reset_req_in8  (1'b0),                                      // (terminated)
		.reset_in9      (1'b0),                                      // (terminated)
		.reset_req_in9  (1'b0),                                      // (terminated)
		.reset_in10     (1'b0),                                      // (terminated)
		.reset_req_in10 (1'b0),                                      // (terminated)
		.reset_in11     (1'b0),                                      // (terminated)
		.reset_req_in11 (1'b0),                                      // (terminated)
		.reset_in12     (1'b0),                                      // (terminated)
		.reset_req_in12 (1'b0),                                      // (terminated)
		.reset_in13     (1'b0),                                      // (terminated)
		.reset_req_in13 (1'b0),                                      // (terminated)
		.reset_in14     (1'b0),                                      // (terminated)
		.reset_req_in14 (1'b0),                                      // (terminated)
		.reset_in15     (1'b0),                                      // (terminated)
		.reset_req_in15 (1'b0)                                       // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
