// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Tue Jun 27 20:09:09 2023"

module RansacNios(
	CLOCK_50,
	KEY,
	receiver_data,
	sender_data
);


input wire	CLOCK_50;
input wire	[0:0] KEY;
input wire	[31:0] receiver_data;
output wire	[31:0] sender_data;






SistemaEmbarcadoRansac	b2v_inst(
	.clk_clk(CLOCK_50),
	.reset_reset_n(KEY),
	.receiver_data_export(receiver_data),
	.sender_data_export(sender_data));


endmodule
