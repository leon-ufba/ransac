
module SistemaEmbarcado (
	clk_clk,
	reset_reset_n,
	medidordesempenho_readdata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[31:0]	medidordesempenho_readdata;
endmodule
