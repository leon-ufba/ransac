// SistemaEmbarcado_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcado_tb (
	);

	wire         sistemaembarcado_inst_clk_bfm_clk_clk;                    // SistemaEmbarcado_inst_clk_bfm:clk -> [SistemaEmbarcado_inst:clk_clk, SistemaEmbarcado_inst_medidordesempenho_conduit_bfm:clk, SistemaEmbarcado_inst_reset_bfm:clk]
	wire  [31:0] sistemaembarcado_inst_medidordesempenho_conduit_readdata; // SistemaEmbarcado_inst:medidordesempenho_conduit_readdata -> SistemaEmbarcado_inst_medidordesempenho_conduit_bfm:sig_readdata
	wire         sistemaembarcado_inst_reset_bfm_reset_reset;              // SistemaEmbarcado_inst_reset_bfm:reset -> [SistemaEmbarcado_inst:reset_reset_n, SistemaEmbarcado_inst_medidordesempenho_conduit_bfm:reset]

	SistemaEmbarcado sistemaembarcado_inst (
		.clk_clk                            (sistemaembarcado_inst_clk_bfm_clk_clk),                    //                       clk.clk
		.medidordesempenho_conduit_readdata (sistemaembarcado_inst_medidordesempenho_conduit_readdata), // medidordesempenho_conduit.readdata
		.reset_reset_n                      (sistemaembarcado_inst_reset_bfm_reset_reset)               //                     reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sistemaembarcado_inst_clk_bfm (
		.clk (sistemaembarcado_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm sistemaembarcado_inst_medidordesempenho_conduit_bfm (
		.clk          (sistemaembarcado_inst_clk_bfm_clk_clk),                    //     clk.clk
		.reset        (~sistemaembarcado_inst_reset_bfm_reset_reset),             //   reset.reset
		.sig_readdata (sistemaembarcado_inst_medidordesempenho_conduit_readdata)  // conduit.readdata
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sistemaembarcado_inst_reset_bfm (
		.reset (sistemaembarcado_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sistemaembarcado_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
