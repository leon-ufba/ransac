
module RANSAC_NIOS (
	clk_clk,
	reset_reset_n,
	medidordesempenho_conduit_readdata);	

	input		clk_clk;
	input		reset_reset_n;
	output	[31:0]	medidordesempenho_conduit_readdata;
endmodule
