// SistemaEmbarcado_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcado_tb (
	);

	wire    sistemaembarcado_inst_clk_bfm_clk_clk;       // SistemaEmbarcado_inst_clk_bfm:clk -> [SistemaEmbarcado_inst:clk_clk, SistemaEmbarcado_inst_reset_bfm:clk]
	wire    sistemaembarcado_inst_reset_bfm_reset_reset; // SistemaEmbarcado_inst_reset_bfm:reset -> SistemaEmbarcado_inst:reset_reset_n

	SistemaEmbarcado sistemaembarcado_inst (
		.clk_clk       (sistemaembarcado_inst_clk_bfm_clk_clk),       //   clk.clk
		.reset_reset_n (sistemaembarcado_inst_reset_bfm_reset_reset)  // reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) sistemaembarcado_inst_clk_bfm (
		.clk (sistemaembarcado_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) sistemaembarcado_inst_reset_bfm (
		.reset (sistemaembarcado_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (sistemaembarcado_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
