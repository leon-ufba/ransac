// SistemaEmbarcado.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module SistemaEmbarcado (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         processador_custom_instruction_master_readra;                                      // Processador:D_ci_readra -> Processador_custom_instruction_master_translator:ci_slave_readra
	wire   [4:0] processador_custom_instruction_master_a;                                           // Processador:D_ci_a -> Processador_custom_instruction_master_translator:ci_slave_a
	wire   [4:0] processador_custom_instruction_master_b;                                           // Processador:D_ci_b -> Processador_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] processador_custom_instruction_master_c;                                           // Processador:D_ci_c -> Processador_custom_instruction_master_translator:ci_slave_c
	wire         processador_custom_instruction_master_readrb;                                      // Processador:D_ci_readrb -> Processador_custom_instruction_master_translator:ci_slave_readrb
	wire         processador_custom_instruction_master_clk;                                         // Processador:E_ci_multi_clock -> Processador_custom_instruction_master_translator:ci_slave_multi_clk
	wire  [31:0] processador_custom_instruction_master_ipending;                                    // Processador:W_ci_ipending -> Processador_custom_instruction_master_translator:ci_slave_ipending
	wire         processador_custom_instruction_master_start;                                       // Processador:E_ci_multi_start -> Processador_custom_instruction_master_translator:ci_slave_multi_start
	wire         processador_custom_instruction_master_reset_req;                                   // Processador:E_ci_multi_reset_req -> Processador_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire         processador_custom_instruction_master_done;                                        // Processador_custom_instruction_master_translator:ci_slave_multi_done -> Processador:E_ci_multi_done
	wire   [7:0] processador_custom_instruction_master_n;                                           // Processador:D_ci_n -> Processador_custom_instruction_master_translator:ci_slave_n
	wire  [31:0] processador_custom_instruction_master_result;                                      // Processador_custom_instruction_master_translator:ci_slave_result -> Processador:E_ci_result
	wire         processador_custom_instruction_master_estatus;                                     // Processador:W_ci_estatus -> Processador_custom_instruction_master_translator:ci_slave_estatus
	wire         processador_custom_instruction_master_clk_en;                                      // Processador:E_ci_multi_clk_en -> Processador_custom_instruction_master_translator:ci_slave_multi_clken
	wire  [31:0] processador_custom_instruction_master_datab;                                       // Processador:E_ci_datab -> Processador_custom_instruction_master_translator:ci_slave_datab
	wire  [31:0] processador_custom_instruction_master_dataa;                                       // Processador:E_ci_dataa -> Processador_custom_instruction_master_translator:ci_slave_dataa
	wire         processador_custom_instruction_master_reset;                                       // Processador:E_ci_multi_reset -> Processador_custom_instruction_master_translator:ci_slave_multi_reset
	wire         processador_custom_instruction_master_writerc;                                     // Processador:D_ci_writerc -> Processador_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] processador_custom_instruction_master_translator_comb_ci_master_result;            // Processador_custom_instruction_master_comb_xconnect:ci_slave_result -> Processador_custom_instruction_master_translator:comb_ci_master_result
	wire         processador_custom_instruction_master_translator_comb_ci_master_readra;            // Processador_custom_instruction_master_translator:comb_ci_master_readra -> Processador_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [4:0] processador_custom_instruction_master_translator_comb_ci_master_a;                 // Processador_custom_instruction_master_translator:comb_ci_master_a -> Processador_custom_instruction_master_comb_xconnect:ci_slave_a
	wire   [4:0] processador_custom_instruction_master_translator_comb_ci_master_b;                 // Processador_custom_instruction_master_translator:comb_ci_master_b -> Processador_custom_instruction_master_comb_xconnect:ci_slave_b
	wire         processador_custom_instruction_master_translator_comb_ci_master_readrb;            // Processador_custom_instruction_master_translator:comb_ci_master_readrb -> Processador_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire   [4:0] processador_custom_instruction_master_translator_comb_ci_master_c;                 // Processador_custom_instruction_master_translator:comb_ci_master_c -> Processador_custom_instruction_master_comb_xconnect:ci_slave_c
	wire         processador_custom_instruction_master_translator_comb_ci_master_estatus;           // Processador_custom_instruction_master_translator:comb_ci_master_estatus -> Processador_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] processador_custom_instruction_master_translator_comb_ci_master_ipending;          // Processador_custom_instruction_master_translator:comb_ci_master_ipending -> Processador_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire  [31:0] processador_custom_instruction_master_translator_comb_ci_master_datab;             // Processador_custom_instruction_master_translator:comb_ci_master_datab -> Processador_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] processador_custom_instruction_master_translator_comb_ci_master_dataa;             // Processador_custom_instruction_master_translator:comb_ci_master_dataa -> Processador_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire         processador_custom_instruction_master_translator_comb_ci_master_writerc;           // Processador_custom_instruction_master_translator:comb_ci_master_writerc -> Processador_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire   [7:0] processador_custom_instruction_master_translator_comb_ci_master_n;                 // Processador_custom_instruction_master_translator:comb_ci_master_n -> Processador_custom_instruction_master_comb_xconnect:ci_slave_n
	wire  [31:0] processador_custom_instruction_master_comb_xconnect_ci_master0_result;             // Processador_custom_instruction_master_comb_slave_translator0:ci_slave_result -> Processador_custom_instruction_master_comb_xconnect:ci_master0_result
	wire         processador_custom_instruction_master_comb_xconnect_ci_master0_readra;             // Processador_custom_instruction_master_comb_xconnect:ci_master0_readra -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [4:0] processador_custom_instruction_master_comb_xconnect_ci_master0_a;                  // Processador_custom_instruction_master_comb_xconnect:ci_master0_a -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire   [4:0] processador_custom_instruction_master_comb_xconnect_ci_master0_b;                  // Processador_custom_instruction_master_comb_xconnect:ci_master0_b -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire         processador_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // Processador_custom_instruction_master_comb_xconnect:ci_master0_readrb -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire   [4:0] processador_custom_instruction_master_comb_xconnect_ci_master0_c;                  // Processador_custom_instruction_master_comb_xconnect:ci_master0_c -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire         processador_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // Processador_custom_instruction_master_comb_xconnect:ci_master0_estatus -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] processador_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // Processador_custom_instruction_master_comb_xconnect:ci_master0_ipending -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire  [31:0] processador_custom_instruction_master_comb_xconnect_ci_master0_datab;              // Processador_custom_instruction_master_comb_xconnect:ci_master0_datab -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] processador_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // Processador_custom_instruction_master_comb_xconnect:ci_master0_dataa -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire         processador_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // Processador_custom_instruction_master_comb_xconnect:ci_master0_writerc -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire   [7:0] processador_custom_instruction_master_comb_xconnect_ci_master0_n;                  // Processador_custom_instruction_master_comb_xconnect:ci_master0_n -> Processador_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire  [31:0] processador_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios_custom_instr_floating_point_2_0:s1_result -> Processador_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] processador_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // Processador_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] processador_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // Processador_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] processador_custom_instruction_master_comb_slave_translator0_ci_master_n;          // Processador_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire         processador_custom_instruction_master_translator_multi_ci_master_readra;           // Processador_custom_instruction_master_translator:multi_ci_master_readra -> Processador_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire   [4:0] processador_custom_instruction_master_translator_multi_ci_master_a;                // Processador_custom_instruction_master_translator:multi_ci_master_a -> Processador_custom_instruction_master_multi_xconnect:ci_slave_a
	wire   [4:0] processador_custom_instruction_master_translator_multi_ci_master_b;                // Processador_custom_instruction_master_translator:multi_ci_master_b -> Processador_custom_instruction_master_multi_xconnect:ci_slave_b
	wire         processador_custom_instruction_master_translator_multi_ci_master_clk;              // Processador_custom_instruction_master_translator:multi_ci_master_clk -> Processador_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         processador_custom_instruction_master_translator_multi_ci_master_readrb;           // Processador_custom_instruction_master_translator:multi_ci_master_readrb -> Processador_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire   [4:0] processador_custom_instruction_master_translator_multi_ci_master_c;                // Processador_custom_instruction_master_translator:multi_ci_master_c -> Processador_custom_instruction_master_multi_xconnect:ci_slave_c
	wire         processador_custom_instruction_master_translator_multi_ci_master_start;            // Processador_custom_instruction_master_translator:multi_ci_master_start -> Processador_custom_instruction_master_multi_xconnect:ci_slave_start
	wire         processador_custom_instruction_master_translator_multi_ci_master_reset_req;        // Processador_custom_instruction_master_translator:multi_ci_master_reset_req -> Processador_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         processador_custom_instruction_master_translator_multi_ci_master_done;             // Processador_custom_instruction_master_multi_xconnect:ci_slave_done -> Processador_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] processador_custom_instruction_master_translator_multi_ci_master_n;                // Processador_custom_instruction_master_translator:multi_ci_master_n -> Processador_custom_instruction_master_multi_xconnect:ci_slave_n
	wire  [31:0] processador_custom_instruction_master_translator_multi_ci_master_result;           // Processador_custom_instruction_master_multi_xconnect:ci_slave_result -> Processador_custom_instruction_master_translator:multi_ci_master_result
	wire         processador_custom_instruction_master_translator_multi_ci_master_clk_en;           // Processador_custom_instruction_master_translator:multi_ci_master_clken -> Processador_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire  [31:0] processador_custom_instruction_master_translator_multi_ci_master_datab;            // Processador_custom_instruction_master_translator:multi_ci_master_datab -> Processador_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire  [31:0] processador_custom_instruction_master_translator_multi_ci_master_dataa;            // Processador_custom_instruction_master_translator:multi_ci_master_dataa -> Processador_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         processador_custom_instruction_master_translator_multi_ci_master_reset;            // Processador_custom_instruction_master_translator:multi_ci_master_reset -> Processador_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire         processador_custom_instruction_master_translator_multi_ci_master_writerc;          // Processador_custom_instruction_master_translator:multi_ci_master_writerc -> Processador_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_readra;            // Processador_custom_instruction_master_multi_xconnect:ci_master0_readra -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire   [4:0] processador_custom_instruction_master_multi_xconnect_ci_master0_a;                 // Processador_custom_instruction_master_multi_xconnect:ci_master0_a -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [4:0] processador_custom_instruction_master_multi_xconnect_ci_master0_b;                 // Processador_custom_instruction_master_multi_xconnect:ci_master0_b -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // Processador_custom_instruction_master_multi_xconnect:ci_master0_readrb -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire   [4:0] processador_custom_instruction_master_multi_xconnect_ci_master0_c;                 // Processador_custom_instruction_master_multi_xconnect:ci_master0_c -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_clk;               // Processador_custom_instruction_master_multi_xconnect:ci_master0_clk -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire  [31:0] processador_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // Processador_custom_instruction_master_multi_xconnect:ci_master0_ipending -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_start;             // Processador_custom_instruction_master_multi_xconnect:ci_master0_start -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // Processador_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_done;              // Processador_custom_instruction_master_multi_slave_translator0:ci_slave_done -> Processador_custom_instruction_master_multi_xconnect:ci_master0_done
	wire   [7:0] processador_custom_instruction_master_multi_xconnect_ci_master0_n;                 // Processador_custom_instruction_master_multi_xconnect:ci_master0_n -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire  [31:0] processador_custom_instruction_master_multi_xconnect_ci_master0_result;            // Processador_custom_instruction_master_multi_slave_translator0:ci_slave_result -> Processador_custom_instruction_master_multi_xconnect:ci_master0_result
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // Processador_custom_instruction_master_multi_xconnect:ci_master0_estatus -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // Processador_custom_instruction_master_multi_xconnect:ci_master0_clken -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire  [31:0] processador_custom_instruction_master_multi_xconnect_ci_master0_datab;             // Processador_custom_instruction_master_multi_xconnect:ci_master0_datab -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire  [31:0] processador_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // Processador_custom_instruction_master_multi_xconnect:ci_master0_dataa -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_reset;             // Processador_custom_instruction_master_multi_xconnect:ci_master0_reset -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire         processador_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // Processador_custom_instruction_master_multi_xconnect:ci_master0_writerc -> Processador_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] processador_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios_custom_instr_floating_point_2_0:s2_result -> Processador_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // Processador_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // Processador_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire  [31:0] processador_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // Processador_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire  [31:0] processador_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // Processador_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_start;     // Processador_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // Processador_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // Processador_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         processador_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios_custom_instr_floating_point_2_0:s2_done -> Processador_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire   [2:0] processador_custom_instruction_master_multi_slave_translator0_ci_master_n;         // Processador_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire  [31:0] processador_data_master_readdata;                                                  // mm_interconnect_0:Processador_data_master_readdata -> Processador:d_readdata
	wire         processador_data_master_waitrequest;                                               // mm_interconnect_0:Processador_data_master_waitrequest -> Processador:d_waitrequest
	wire         processador_data_master_debugaccess;                                               // Processador:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:Processador_data_master_debugaccess
	wire  [18:0] processador_data_master_address;                                                   // Processador:d_address -> mm_interconnect_0:Processador_data_master_address
	wire   [3:0] processador_data_master_byteenable;                                                // Processador:d_byteenable -> mm_interconnect_0:Processador_data_master_byteenable
	wire         processador_data_master_read;                                                      // Processador:d_read -> mm_interconnect_0:Processador_data_master_read
	wire         processador_data_master_write;                                                     // Processador:d_write -> mm_interconnect_0:Processador_data_master_write
	wire  [31:0] processador_data_master_writedata;                                                 // Processador:d_writedata -> mm_interconnect_0:Processador_data_master_writedata
	wire  [31:0] processador_instruction_master_readdata;                                           // mm_interconnect_0:Processador_instruction_master_readdata -> Processador:i_readdata
	wire         processador_instruction_master_waitrequest;                                        // mm_interconnect_0:Processador_instruction_master_waitrequest -> Processador:i_waitrequest
	wire  [18:0] processador_instruction_master_address;                                            // Processador:i_address -> mm_interconnect_0:Processador_instruction_master_address
	wire         processador_instruction_master_read;                                               // Processador:i_read -> mm_interconnect_0:Processador_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_processador_debug_mem_slave_readdata;                            // Processador:debug_mem_slave_readdata -> mm_interconnect_0:Processador_debug_mem_slave_readdata
	wire         mm_interconnect_0_processador_debug_mem_slave_waitrequest;                         // Processador:debug_mem_slave_waitrequest -> mm_interconnect_0:Processador_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_processador_debug_mem_slave_debugaccess;                         // mm_interconnect_0:Processador_debug_mem_slave_debugaccess -> Processador:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_processador_debug_mem_slave_address;                             // mm_interconnect_0:Processador_debug_mem_slave_address -> Processador:debug_mem_slave_address
	wire         mm_interconnect_0_processador_debug_mem_slave_read;                                // mm_interconnect_0:Processador_debug_mem_slave_read -> Processador:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_processador_debug_mem_slave_byteenable;                          // mm_interconnect_0:Processador_debug_mem_slave_byteenable -> Processador:debug_mem_slave_byteenable
	wire         mm_interconnect_0_processador_debug_mem_slave_write;                               // mm_interconnect_0:Processador_debug_mem_slave_write -> Processador:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_processador_debug_mem_slave_writedata;                           // mm_interconnect_0:Processador_debug_mem_slave_writedata -> Processador:debug_mem_slave_writedata
	wire         mm_interconnect_0_memoriaprograma_s1_chipselect;                                   // mm_interconnect_0:MemoriaPrograma_s1_chipselect -> MemoriaPrograma:chipselect
	wire  [31:0] mm_interconnect_0_memoriaprograma_s1_readdata;                                     // MemoriaPrograma:readdata -> mm_interconnect_0:MemoriaPrograma_s1_readdata
	wire  [14:0] mm_interconnect_0_memoriaprograma_s1_address;                                      // mm_interconnect_0:MemoriaPrograma_s1_address -> MemoriaPrograma:address
	wire   [3:0] mm_interconnect_0_memoriaprograma_s1_byteenable;                                   // mm_interconnect_0:MemoriaPrograma_s1_byteenable -> MemoriaPrograma:byteenable
	wire         mm_interconnect_0_memoriaprograma_s1_write;                                        // mm_interconnect_0:MemoriaPrograma_s1_write -> MemoriaPrograma:write
	wire  [31:0] mm_interconnect_0_memoriaprograma_s1_writedata;                                    // mm_interconnect_0:MemoriaPrograma_s1_writedata -> MemoriaPrograma:writedata
	wire         mm_interconnect_0_memoriaprograma_s1_clken;                                        // mm_interconnect_0:MemoriaPrograma_s1_clken -> MemoriaPrograma:clken
	wire         mm_interconnect_0_memoriadados_s1_chipselect;                                      // mm_interconnect_0:MemoriaDados_s1_chipselect -> MemoriaDados:chipselect
	wire  [31:0] mm_interconnect_0_memoriadados_s1_readdata;                                        // MemoriaDados:readdata -> mm_interconnect_0:MemoriaDados_s1_readdata
	wire  [13:0] mm_interconnect_0_memoriadados_s1_address;                                         // mm_interconnect_0:MemoriaDados_s1_address -> MemoriaDados:address
	wire   [3:0] mm_interconnect_0_memoriadados_s1_byteenable;                                      // mm_interconnect_0:MemoriaDados_s1_byteenable -> MemoriaDados:byteenable
	wire         mm_interconnect_0_memoriadados_s1_write;                                           // mm_interconnect_0:MemoriaDados_s1_write -> MemoriaDados:write
	wire  [31:0] mm_interconnect_0_memoriadados_s1_writedata;                                       // mm_interconnect_0:MemoriaDados_s1_writedata -> MemoriaDados:writedata
	wire         mm_interconnect_0_memoriadados_s1_clken;                                           // mm_interconnect_0:MemoriaDados_s1_clken -> MemoriaDados:clken
	wire         irq_mapper_receiver0_irq;                                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] processador_irq_irq;                                                               // irq_mapper:sender_irq -> Processador:irq
	wire         rst_controller_reset_out_reset;                                                    // rst_controller:reset_out -> [MemoriaDados:reset, MemoriaPrograma:reset, Processador:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:Processador_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                                // rst_controller:reset_req -> [MemoriaDados:reset_req, MemoriaPrograma:reset_req, Processador:reset_req, rst_translator:reset_req_in]
	wire         processador_debug_reset_request_reset;                                             // Processador:debug_reset_request -> rst_controller:reset_in1

	SistemaEmbarcado_MemoriaDados memoriadados (
		.clk        (clk_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_memoriadados_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoriadados_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoriadados_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoriadados_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoriadados_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoriadados_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoriadados_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze     (1'b0)                                          // (terminated)
	);

	SistemaEmbarcado_MemoriaPrograma memoriaprograma (
		.clk        (clk_clk),                                         //   clk1.clk
		.address    (mm_interconnect_0_memoriaprograma_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_memoriaprograma_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_memoriaprograma_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_memoriaprograma_s1_write),      //       .write
		.readdata   (mm_interconnect_0_memoriaprograma_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_memoriaprograma_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_memoriaprograma_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),              //       .reset_req
		.freeze     (1'b0)                                             // (terminated)
	);

	SistemaEmbarcado_Processador processador (
		.clk                                 (clk_clk),                                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                           //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                           (processador_data_master_address),                           //               data_master.address
		.d_byteenable                        (processador_data_master_byteenable),                        //                          .byteenable
		.d_read                              (processador_data_master_read),                              //                          .read
		.d_readdata                          (processador_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (processador_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (processador_data_master_write),                             //                          .write
		.d_writedata                         (processador_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (processador_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (processador_instruction_master_address),                    //        instruction_master.address
		.i_read                              (processador_instruction_master_read),                       //                          .read
		.i_readdata                          (processador_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (processador_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (processador_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (processador_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_processador_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_processador_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_processador_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_processador_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_processador_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_processador_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_processador_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_processador_debug_mem_slave_writedata),   //                          .writedata
		.E_ci_multi_done                     (processador_custom_instruction_master_done),                // custom_instruction_master.done
		.E_ci_multi_clk_en                   (processador_custom_instruction_master_clk_en),              //                          .clk_en
		.E_ci_multi_start                    (processador_custom_instruction_master_start),               //                          .start
		.E_ci_result                         (processador_custom_instruction_master_result),              //                          .result
		.D_ci_a                              (processador_custom_instruction_master_a),                   //                          .a
		.D_ci_b                              (processador_custom_instruction_master_b),                   //                          .b
		.D_ci_c                              (processador_custom_instruction_master_c),                   //                          .c
		.D_ci_n                              (processador_custom_instruction_master_n),                   //                          .n
		.D_ci_readra                         (processador_custom_instruction_master_readra),              //                          .readra
		.D_ci_readrb                         (processador_custom_instruction_master_readrb),              //                          .readrb
		.D_ci_writerc                        (processador_custom_instruction_master_writerc),             //                          .writerc
		.E_ci_dataa                          (processador_custom_instruction_master_dataa),               //                          .dataa
		.E_ci_datab                          (processador_custom_instruction_master_datab),               //                          .datab
		.E_ci_multi_clock                    (processador_custom_instruction_master_clk),                 //                          .clk
		.E_ci_multi_reset                    (processador_custom_instruction_master_reset),               //                          .reset
		.E_ci_multi_reset_req                (processador_custom_instruction_master_reset_req),           //                          .reset_req
		.W_ci_estatus                        (processador_custom_instruction_master_estatus),             //                          .estatus
		.W_ci_ipending                       (processador_custom_instruction_master_ipending)             //                          .ipending
	);

	SistemaEmbarcado_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	SistemaEmbarcado_nios_custom_instr_floating_point_2_0 #(
		.arithmetic_present (1),
		.root_present       (0),
		.conversion_present (1),
		.comparison_present (1)
	) nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (processador_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (processador_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (processador_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (processador_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (processador_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (processador_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (processador_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (processador_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (processador_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (processador_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (processador_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (processador_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (processador_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (processador_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (1)
	) processador_custom_instruction_master_translator (
		.ci_slave_dataa            (processador_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (processador_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (processador_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (processador_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (processador_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (processador_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (processador_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (processador_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (processador_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (processador_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (processador_custom_instruction_master_ipending),                             //                .ipending
		.ci_slave_estatus          (processador_custom_instruction_master_estatus),                              //                .estatus
		.ci_slave_multi_clk        (processador_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (processador_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (processador_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (processador_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (processador_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (processador_custom_instruction_master_done),                                 //                .done
		.comb_ci_master_dataa      (processador_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (processador_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (processador_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (processador_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (processador_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (processador_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (processador_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (processador_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (processador_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (processador_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (processador_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (processador_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (processador_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (processador_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (processador_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (processador_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (processador_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (processador_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (processador_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (processador_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (processador_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (processador_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (processador_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (processador_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (processador_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (processador_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (processador_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (processador_custom_instruction_master_translator_multi_ci_master_c),         //                .c
		.ci_slave_multi_dataa      (32'b00000000000000000000000000000000),                                       //     (terminated)
		.ci_slave_multi_datab      (32'b00000000000000000000000000000000),                                       //     (terminated)
		.ci_slave_multi_result     (),                                                                           //     (terminated)
		.ci_slave_multi_n          (8'b00000000),                                                                //     (terminated)
		.ci_slave_multi_readra     (1'b0),                                                                       //     (terminated)
		.ci_slave_multi_readrb     (1'b0),                                                                       //     (terminated)
		.ci_slave_multi_writerc    (1'b0),                                                                       //     (terminated)
		.ci_slave_multi_a          (5'b00000),                                                                   //     (terminated)
		.ci_slave_multi_b          (5'b00000),                                                                   //     (terminated)
		.ci_slave_multi_c          (5'b00000)                                                                    //     (terminated)
	);

	SistemaEmbarcado_Processador_custom_instruction_master_comb_xconnect processador_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (processador_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (processador_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (processador_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (processador_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (processador_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (processador_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (processador_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (processador_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (processador_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (processador_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (processador_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (processador_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (processador_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (processador_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (processador_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (processador_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (processador_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (processador_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (processador_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (processador_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (processador_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (processador_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (processador_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (processador_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) processador_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (processador_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (processador_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (processador_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (processador_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (processador_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (processador_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (processador_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (processador_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (processador_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (processador_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (processador_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (processador_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (processador_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (processador_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (processador_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (processador_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                              // (terminated)
		.ci_master_readrb    (),                                                                              // (terminated)
		.ci_master_writerc   (),                                                                              // (terminated)
		.ci_master_a         (),                                                                              // (terminated)
		.ci_master_b         (),                                                                              // (terminated)
		.ci_master_c         (),                                                                              // (terminated)
		.ci_master_ipending  (),                                                                              // (terminated)
		.ci_master_estatus   (),                                                                              // (terminated)
		.ci_master_clk       (),                                                                              // (terminated)
		.ci_master_clken     (),                                                                              // (terminated)
		.ci_master_reset_req (),                                                                              // (terminated)
		.ci_master_reset     (),                                                                              // (terminated)
		.ci_master_start     (),                                                                              // (terminated)
		.ci_master_done      (1'b0),                                                                          // (terminated)
		.ci_slave_clk        (1'b0),                                                                          // (terminated)
		.ci_slave_clken      (1'b0),                                                                          // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                          // (terminated)
		.ci_slave_reset      (1'b0),                                                                          // (terminated)
		.ci_slave_start      (1'b0),                                                                          // (terminated)
		.ci_slave_done       ()                                                                               // (terminated)
	);

	SistemaEmbarcado_Processador_custom_instruction_master_multi_xconnect processador_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (processador_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (processador_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (processador_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (processador_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (processador_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (processador_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (processador_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (processador_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (processador_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (processador_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                           //           .ipending
		.ci_slave_estatus     (),                                                                           //           .estatus
		.ci_slave_clk         (processador_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (processador_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (processador_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (processador_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (processador_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (processador_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (processador_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (processador_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (processador_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (processador_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (processador_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (processador_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (processador_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (processador_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (processador_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (processador_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (processador_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (processador_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (processador_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (processador_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (processador_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (processador_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (processador_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (processador_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) processador_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (processador_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (processador_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (processador_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (processador_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (processador_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (processador_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (processador_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (processador_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (processador_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (processador_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (processador_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (processador_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (processador_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (processador_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (processador_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (processador_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (processador_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (processador_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (processador_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (processador_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (processador_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (processador_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (processador_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (processador_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (processador_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (processador_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (processador_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (processador_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                                  // (terminated)
		.ci_master_readrb    (),                                                                                  // (terminated)
		.ci_master_writerc   (),                                                                                  // (terminated)
		.ci_master_a         (),                                                                                  // (terminated)
		.ci_master_b         (),                                                                                  // (terminated)
		.ci_master_c         (),                                                                                  // (terminated)
		.ci_master_ipending  (),                                                                                  // (terminated)
		.ci_master_estatus   ()                                                                                   // (terminated)
	);

	SistemaEmbarcado_mm_interconnect_0 mm_interconnect_0 (
		.clock_clk_clk                                 (clk_clk),                                                   //                               clock_clk.clk
		.Processador_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // Processador_reset_reset_bridge_in_reset.reset
		.Processador_data_master_address               (processador_data_master_address),                           //                 Processador_data_master.address
		.Processador_data_master_waitrequest           (processador_data_master_waitrequest),                       //                                        .waitrequest
		.Processador_data_master_byteenable            (processador_data_master_byteenable),                        //                                        .byteenable
		.Processador_data_master_read                  (processador_data_master_read),                              //                                        .read
		.Processador_data_master_readdata              (processador_data_master_readdata),                          //                                        .readdata
		.Processador_data_master_write                 (processador_data_master_write),                             //                                        .write
		.Processador_data_master_writedata             (processador_data_master_writedata),                         //                                        .writedata
		.Processador_data_master_debugaccess           (processador_data_master_debugaccess),                       //                                        .debugaccess
		.Processador_instruction_master_address        (processador_instruction_master_address),                    //          Processador_instruction_master.address
		.Processador_instruction_master_waitrequest    (processador_instruction_master_waitrequest),                //                                        .waitrequest
		.Processador_instruction_master_read           (processador_instruction_master_read),                       //                                        .read
		.Processador_instruction_master_readdata       (processador_instruction_master_readdata),                   //                                        .readdata
		.jtag_uart_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.jtag_uart_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.jtag_uart_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.MemoriaDados_s1_address                       (mm_interconnect_0_memoriadados_s1_address),                 //                         MemoriaDados_s1.address
		.MemoriaDados_s1_write                         (mm_interconnect_0_memoriadados_s1_write),                   //                                        .write
		.MemoriaDados_s1_readdata                      (mm_interconnect_0_memoriadados_s1_readdata),                //                                        .readdata
		.MemoriaDados_s1_writedata                     (mm_interconnect_0_memoriadados_s1_writedata),               //                                        .writedata
		.MemoriaDados_s1_byteenable                    (mm_interconnect_0_memoriadados_s1_byteenable),              //                                        .byteenable
		.MemoriaDados_s1_chipselect                    (mm_interconnect_0_memoriadados_s1_chipselect),              //                                        .chipselect
		.MemoriaDados_s1_clken                         (mm_interconnect_0_memoriadados_s1_clken),                   //                                        .clken
		.MemoriaPrograma_s1_address                    (mm_interconnect_0_memoriaprograma_s1_address),              //                      MemoriaPrograma_s1.address
		.MemoriaPrograma_s1_write                      (mm_interconnect_0_memoriaprograma_s1_write),                //                                        .write
		.MemoriaPrograma_s1_readdata                   (mm_interconnect_0_memoriaprograma_s1_readdata),             //                                        .readdata
		.MemoriaPrograma_s1_writedata                  (mm_interconnect_0_memoriaprograma_s1_writedata),            //                                        .writedata
		.MemoriaPrograma_s1_byteenable                 (mm_interconnect_0_memoriaprograma_s1_byteenable),           //                                        .byteenable
		.MemoriaPrograma_s1_chipselect                 (mm_interconnect_0_memoriaprograma_s1_chipselect),           //                                        .chipselect
		.MemoriaPrograma_s1_clken                      (mm_interconnect_0_memoriaprograma_s1_clken),                //                                        .clken
		.Processador_debug_mem_slave_address           (mm_interconnect_0_processador_debug_mem_slave_address),     //             Processador_debug_mem_slave.address
		.Processador_debug_mem_slave_write             (mm_interconnect_0_processador_debug_mem_slave_write),       //                                        .write
		.Processador_debug_mem_slave_read              (mm_interconnect_0_processador_debug_mem_slave_read),        //                                        .read
		.Processador_debug_mem_slave_readdata          (mm_interconnect_0_processador_debug_mem_slave_readdata),    //                                        .readdata
		.Processador_debug_mem_slave_writedata         (mm_interconnect_0_processador_debug_mem_slave_writedata),   //                                        .writedata
		.Processador_debug_mem_slave_byteenable        (mm_interconnect_0_processador_debug_mem_slave_byteenable),  //                                        .byteenable
		.Processador_debug_mem_slave_waitrequest       (mm_interconnect_0_processador_debug_mem_slave_waitrequest), //                                        .waitrequest
		.Processador_debug_mem_slave_debugaccess       (mm_interconnect_0_processador_debug_mem_slave_debugaccess)  //                                        .debugaccess
	);

	SistemaEmbarcado_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (processador_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                        // reset_in0.reset
		.reset_in1      (processador_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                               //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),    //          .reset_req
		.reset_req_in0  (1'b0),                                  // (terminated)
		.reset_req_in1  (1'b0),                                  // (terminated)
		.reset_in2      (1'b0),                                  // (terminated)
		.reset_req_in2  (1'b0),                                  // (terminated)
		.reset_in3      (1'b0),                                  // (terminated)
		.reset_req_in3  (1'b0),                                  // (terminated)
		.reset_in4      (1'b0),                                  // (terminated)
		.reset_req_in4  (1'b0),                                  // (terminated)
		.reset_in5      (1'b0),                                  // (terminated)
		.reset_req_in5  (1'b0),                                  // (terminated)
		.reset_in6      (1'b0),                                  // (terminated)
		.reset_req_in6  (1'b0),                                  // (terminated)
		.reset_in7      (1'b0),                                  // (terminated)
		.reset_req_in7  (1'b0),                                  // (terminated)
		.reset_in8      (1'b0),                                  // (terminated)
		.reset_req_in8  (1'b0),                                  // (terminated)
		.reset_in9      (1'b0),                                  // (terminated)
		.reset_req_in9  (1'b0),                                  // (terminated)
		.reset_in10     (1'b0),                                  // (terminated)
		.reset_req_in10 (1'b0),                                  // (terminated)
		.reset_in11     (1'b0),                                  // (terminated)
		.reset_req_in11 (1'b0),                                  // (terminated)
		.reset_in12     (1'b0),                                  // (terminated)
		.reset_req_in12 (1'b0),                                  // (terminated)
		.reset_in13     (1'b0),                                  // (terminated)
		.reset_req_in13 (1'b0),                                  // (terminated)
		.reset_in14     (1'b0),                                  // (terminated)
		.reset_req_in14 (1'b0),                                  // (terminated)
		.reset_in15     (1'b0),                                  // (terminated)
		.reset_req_in15 (1'b0)                                   // (terminated)
	);

endmodule
